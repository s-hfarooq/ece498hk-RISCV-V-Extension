
module digitalTimer (
    input logic clk,
    input logic rst
);

endmodule : digitalTimer
