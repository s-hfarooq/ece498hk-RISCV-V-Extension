
module sram (
    input logic clk,
    input logic rst
);

endmodule : sram
