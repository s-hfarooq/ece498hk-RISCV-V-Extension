
module spi (
    input logic clk,
    input logic rst
);

endmodule : spi
