module io_buf (
    input   logic   i,
    output  logic   o
);

buf (o, i);

endmodule