
module uart (
    input logic clk,
    input logic rst
);

endmodule : uart
